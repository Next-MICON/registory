module hardware (
    // Left side
    inout pin1,
    inout pin2,
    inout pin3,
    inout pin4,
    inout pin5,
    inout pin6,
    inout pin7,
    inout pin8,
    inout pin9,
    inout pin10,
    inout pin11,
    inout pin12,
    inout pin13,

    // Right side
    inout pin14,
    inout pin15,
    inout pin16,
    inout pin17,
    inout pin18,
    inout pin19,
    inout pin20,
    inout pin21,
    inout pin22,
    inout pin23,
    inout pin24,

    // Bottom
    inout pin25,
    inout pin26,
    inout pin27,
    inout pin28,
    inout pin29,
    inout pin30,
    inout pin31,

    // SPI Flash
    inout flash_csb,
    inout flash_clk,
    inout flash_io0,
    inout flash_io1,
    inout flash_io2,
    inout flash_io3,

    // LED
    inout led,

    // USB
    inout usb_pu,
    inout usb_p,
    inout usb_n,

    // Clock
    input clk_16MHz
);

  /* iobuffer */
  /* end */

  ///////////////////////////////////
  // Clock & Reset

  por por (
      .clk(clk),
      .resetn(resetn)
  );
  wire clk = clk_16MHz;
  wire resetn;

  ///////////////////////////////////
  // Parameters

  parameter integer MEM_WORDS = 2048;
  parameter [31:0] STACKADDR = (4 * MEM_WORDS);  // end of memory
  parameter [31:0] PROGADDR_RESET = 32'h0005_0000;  // 1 MB into flash
  parameter [31:0] PROGADDR_IRQ = 32'h0005_0010;  // 1 MB into flash

  /* parameters */
  /* end */

  ///////////////////////////////////
  // Interrupts Request

  reg [31:0] irq;
  always @* begin
    if (!resetn) irq <= 0;
    else begin
      irq = 0;
      /* irq */
      irq[5] = pin11;
      /* end */
    end
  end

  ///////////////////////////////////
  // CPU

  picorv32 #(
      .STACKADDR(STACKADDR),
      .PROGADDR_RESET(PROGADDR_RESET),
      .PROGADDR_IRQ(PROGADDR_IRQ),
      .BARREL_SHIFTER(1),
      .COMPRESSED_ISA(1),
      .ENABLE_MUL(1),
      .ENABLE_DIV(1),
      .ENABLE_IRQ(1),
      .ENABLE_IRQ_QREGS(1)
  ) cpu (
      .clk      (clk),
      .resetn   (resetn),
      .mem_valid(mem_valid),
      .mem_ready(mem_ready),
      .mem_addr (mem_addr),
      .mem_wdata(mem_wdata),
      .mem_wstrb(mem_wstrb),
      .mem_rdata(mem_rdata),
      .irq      (irq)
  );

  ///////////////////////////////////
  // Memory map interface

  wire mem_valid;
  wire mem_ready;
  wire [3:0] mem_wstrb;
  wire [31:0] mem_addr;
  wire [31:0] mem_wdata;
  wire [31:0] mem_rdata;
  assign mem_ready = |{ram_ready, rom_ready, rom_cfg_ready
      /* mem_ready */
      /* end */};
  assign mem_rdata = ram_ready ? ram_rdata : rom_ready ? rom_rdata : rom_cfg_ready ? rom_cfg_rdata
      /* mem_rdata */
      /* end */ : 32'b0;

  ///////////////////////////////////
  // Modules

  ram #(
      .WORDS(MEM_WORDS)
  ) ram (
      .clk(clk),
      .resetn(resetn),
      .valid(ram_valid),
      .ready(ram_ready),
      .wstrb(ram_valid ? mem_wstrb : 4'b0),
      .addr(mem_addr),
      .wdata(mem_wdata),
      .rdata(ram_rdata)
  );
  wire ram_sel = mem_addr[31:14] == 19'h0;
  wire ram_valid = mem_valid && ram_sel;
  wire ram_ready;
  wire [31:0] ram_rdata;

  spirom rom (
      .clk(clk),
      .resetn(resetn),
      .valid(rom_valid),
      .ready(rom_ready),
      .wstrb(rom_valid ? mem_wstrb : 4'b0),
      .addr (mem_addr),
      .wdata(mem_wdata),
      .rdata(rom_rdata),
      .cfg_valid(rom_cfg_valid),
      .cfg_ready(rom_cfg_ready),
      .cfg_wstrb(rom_cfg_valid ? mem_wstrb : 4'b0),
      .cfg_addr (mem_addr),
      .cfg_wdata(mem_wdata),
      .cfg_rdata(rom_cfg_rdata),
      .flash_io0_iosel(flash_io0_iosel),
      .flash_io0_in   (flash_io0_in),
      .flash_io0_out  (flash_io0_out),
      .flash_io1_iosel(flash_io1_iosel),
      .flash_io1_in   (flash_io1_in),
      .flash_io1_out  (flash_io1_out),
      .flash_io2_iosel(flash_io2_iosel),
      .flash_io2_in   (flash_io2_in),
      .flash_io2_out  (flash_io2_out),
      .flash_io3_iosel(flash_io3_iosel),
      .flash_io3_in   (flash_io3_in),
      .flash_io3_out  (flash_io3_out),
      .flash_csb(flash_csb),
      .flash_clk(flash_clk)
  );
  wire rom_sel = (mem_addr[31:20] == 12'h000) && (4'h5 <= mem_addr[19:16]);
  wire rom_valid = mem_valid && rom_sel;
  wire rom_ready;
  wire [31:0] rom_rdata;
  wire rom_cfg_sel = mem_addr[31:24] == 8'h02;
  wire rom_cfg_valid = mem_valid && rom_cfg_sel;
  wire rom_cfg_ready;
  wire [31:0] rom_cfg_rdata;
  wire flash_io0_iosel;
  wire flash_io0_in;
  wire flash_io0_out;
  wire flash_io1_iosel;
  wire flash_io1_in;
  wire flash_io1_out;
  wire flash_io2_iosel;
  wire flash_io2_in;
  wire flash_io2_out;
  wire flash_io3_iosel;
  wire flash_io3_in;
  wire flash_io3_out;
  PortInOut flash_io0_iobuf (
      .pin  (flash_io0),
      .iosel(flash_io0_iosel),
      .out  (flash_io0_in),
      .in   (flash_io0_out)
  );
  PortInOut flash_io1_iobuf (
      .pin  (flash_io1),
      .iosel(flash_io1_iosel),
      .out  (flash_io1_in),
      .in   (flash_io1_out)
  );
  PortInOut flash_io2_iobuf (
      .pin  (flash_io2),
      .iosel(flash_io2_iosel),
      .out  (flash_io2_in),
      .in   (flash_io2_out)
  );
  PortInOut flash_io3_iobuf (
      .pin  (flash_io3),
      .iosel(flash_io3_iosel),
      .out  (flash_io3_in),
      .in   (flash_io3_out)
  );

  /* instances */
  /* end */

endmodule
