module hardware (
    // Left side
    inout pin1,
    inout pin2,
    inout pin3,
    inout pin4,
    inout pin5,
    inout pin6,
    inout pin7,
    inout pin8,
    inout pin9,
    inout pin10,
    inout pin11,
    inout pin12,
    inout pin13,

    // Right side
    inout pin14,
    inout pin15,
    inout pin16,
    inout pin17,
    inout pin18,
    inout pin19,
    inout pin20,
    inout pin21,
    inout pin22,
    inout pin23,
    inout pin24,

    // Bottom
    inout pin25,
    inout pin26,
    inout pin27,
    inout pin28,
    inout pin29,
    inout pin30,
    inout pin31,

    // SPI Flash
    inout flash_csb,
    inout flash_clk,
    inout flash_io0,
    inout flash_io1,
    inout flash_io2,
    inout flash_io3,

    // LED
    inout led,

    // USB
    inout usb_pu,
    inout usb_p,
    inout usb_n,

    // Clock
    input clk_16MHz
);

  /* iobuffer */
In pin2_iobuf(
  .pin(pin2),
  .in(pin2_in)
);
wire pin2_in;
Out pin1_iobuf(
  .pin(pin1),
  .out(serial_tx)
);
InOut pin3_iobuf(
  .pin(pin3),
  .iosel(digital_iosel),
  .out(digital_out),
  .in(pin3_in)
);
wire pin3_in;
Out led_iobuf(
  .pin(led),
  .out(digital_out)
);
In pin11_iobuf(
  .pin(pin11),
  .in(pin11_in)
);
wire pin11_in;
/* end */

  ///////////////////////////////////
  // Wire Deffinitions

  wire clk = clk_16MHz;
  wire resetn;

  ///////////////////////////////////
  // Parameters

  parameter integer MEM_WORDS = 2048;
  parameter [31:0] STACKADDR = (4 * MEM_WORDS);  // end of memory
  parameter [31:0] PROGADDR_RESET = 32'h0005_0000;  // 1 MB into flash
  parameter [31:0] PROGADDR_IRQ = 32'h0005_0010;  // 1 MB into flash

  /* parameters */
  /* end */

  ///////////////////////////////////
  // Interrupts Request

  reg [31:0] irq;
  always @* begin
    if (!resetn) irq <= 0;
    else begin
      irq = 0;
      /* irq */
      irq[3] = pin11_in;
/* end */
    end
  end

  ///////////////////////////////////
  // CPU

  picorv32 #(
      .STACKADDR(STACKADDR),
      .PROGADDR_RESET(PROGADDR_RESET),
      .PROGADDR_IRQ(PROGADDR_IRQ),
      .BARREL_SHIFTER(1),
      .COMPRESSED_ISA(1),
      .ENABLE_MUL(1),
      .ENABLE_DIV(1),
      .ENABLE_IRQ(1),
      .ENABLE_IRQ_QREGS(1)
  ) cpu (
      .clk      (clk),
      .resetn   (resetn),
      .mem_valid(mem_valid),
      .mem_ready(mem_ready),
      .mem_addr (mem_addr),
      .mem_wdata(mem_wdata),
      .mem_wstrb(mem_wstrb),
      .mem_rdata(mem_rdata),
      .irq      (irq)
  );

  ///////////////////////////////////
  // Memory map interface

  wire mem_valid;
  wire mem_ready;
  wire [3:0] mem_wstrb;
  wire [31:0] mem_addr;
  wire [31:0] mem_wdata;
  wire [31:0] mem_rdata;
  assign mem_ready = |{ram_ready, rom_ready, rom_cfg_ready
      /* mem_ready */
, serial_ready, digital_ready
/* end */};
  assign mem_rdata = ram_ready ? ram_rdata : rom_ready ? rom_rdata : rom_cfg_ready ? rom_cfg_rdata
      /* mem_rdata */
: serial_ready ? serial_rdata: digital_ready ? digital_rdata
/* end */ : 32'b0;

  ///////////////////////////////////
  // Modules

  por por (
      .clk(clk),
      .resetn(resetn)
  );

  ram #(
      .WORDS(MEM_WORDS)
  ) ram (
      .clk(clk),
      .resetn(resetn),
      .valid(ram_valid),
      .ready(ram_ready),
      .wstrb(ram_valid ? mem_wstrb : 4'b0),
      .addr(mem_addr),
      .wdata(mem_wdata),
      .rdata(ram_rdata)
  );
  wire ram_sel = mem_addr[31:14] == 19'h0;
  wire ram_valid = mem_valid && ram_sel;
  wire ram_ready;
  wire [31:0] ram_rdata;

  spirom rom (
      .clk(clk),
      .resetn(resetn),
      .valid(rom_valid),
      .ready(rom_ready),
      .wstrb(rom_valid ? mem_wstrb : 4'b0),
      .addr (mem_addr),
      .wdata(mem_wdata),
      .rdata(rom_rdata),
      .cfg_valid(rom_cfg_valid),
      .cfg_ready(rom_cfg_ready),
      .cfg_wstrb(rom_cfg_valid ? mem_wstrb : 4'b0),
      .cfg_addr (mem_addr),
      .cfg_wdata(mem_wdata),
      .cfg_rdata(rom_cfg_rdata),
      .flash_io0_iosel(flash_io0_iosel),
      .flash_io0_in   (flash_io0_in),
      .flash_io0_out  (flash_io0_out),
      .flash_io1_iosel(flash_io1_iosel),
      .flash_io1_in   (flash_io1_in),
      .flash_io1_out  (flash_io1_out),
      .flash_io2_iosel(flash_io2_iosel),
      .flash_io2_in   (flash_io2_in),
      .flash_io2_out  (flash_io2_out),
      .flash_io3_iosel(flash_io3_iosel),
      .flash_io3_in   (flash_io3_in),
      .flash_io3_out  (flash_io3_out),
      .flash_csb(flash_csb),
      .flash_clk(flash_clk)
  );
  wire rom_sel = (mem_addr[31:20] == 12'h000) && (4'h5 <= mem_addr[19:16]);
  wire rom_valid = mem_valid && rom_sel;
  wire rom_ready;
  wire [31:0] rom_rdata;
  wire rom_cfg_sel = mem_addr[31:24] == 8'h02;
  wire rom_cfg_valid = mem_valid && rom_cfg_sel;
  wire rom_cfg_ready;
  wire [31:0] rom_cfg_rdata;
  wire flash_io0_iosel;
  wire flash_io0_in;
  wire flash_io0_out;
  wire flash_io1_iosel;
  wire flash_io1_in;
  wire flash_io1_out;
  wire flash_io2_iosel;
  wire flash_io2_in;
  wire flash_io2_out;
  wire flash_io3_iosel;
  wire flash_io3_in;
  wire flash_io3_out;
  InOut flash_io0_iobuf (
      .pin  (flash_io0),
      .iosel(flash_io0_iosel),
      .in   (flash_io0_in),
      .out  (flash_io0_out)
  );
  InOut flash_io1_iobuf (
      .pin  (flash_io1),
      .iosel(flash_io1_iosel),
      .in   (flash_io1_in),
      .out  (flash_io1_out)
  );
  InOut flash_io2_iobuf (
      .pin  (flash_io2),
      .iosel(flash_io2_iosel),
      .in   (flash_io2_in),
      .out  (flash_io2_out)
  );
  InOut flash_io3_iobuf (
      .pin  (flash_io3),
      .iosel(flash_io3_iosel),
      .in   (flash_io3_in),
      .out  (flash_io3_out)
  );

  /* instances */
Serial serial(
  .clk(clk),
  .resetn(resetn),
  .valid(serial_valid),
  .ready(serial_ready),
  .wstrb(serial_valid ? mem_wstrb : 4'b0),
  .addr(mem_addr),
  .wdata(mem_wdata),
  .rdata(serial_rdata),
  .rx(pin2_in),
  .tx(serial_tx)
);
wire serial_sel = mem_addr[31:24] == 8'h3;
wire serial_valid = mem_valid && serial_sel;
wire serial_ready;
wire [31:0] serial_rdata;
wire serial_tx;

Digital digital(
  .clk(clk),
  .resetn(resetn),
  .valid(digital_valid),
  .ready(digital_ready),
  .wstrb(digital_valid ? mem_wstrb : 4'b0),
  .addr(mem_addr),
  .wdata(mem_wdata),
  .rdata(digital_rdata),
  .iosel(digital_iosel),
  .out(digital_out),
  .in(pin3_in)
);
wire digital_sel = mem_addr[31:24] == 8'h4;
wire digital_valid = mem_valid && digital_sel;
wire digital_ready;
wire [31:0] digital_rdata;
wire digital_iosel;
wire digital_out;
/* end */

endmodule
